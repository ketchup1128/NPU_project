module entry_state #(
    parameters
) (
    input clk, 
    input rst_n, 

    input start,
    input  
    input wr_en, 
);
    
endmodule